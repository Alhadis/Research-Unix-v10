a,b
ab
abcde
alphanum
ARB
ARBNO
binaryop
BREAKX
bstj
cacm
cdr
cstr
DATATYPE
datatype
dequeue
dliteral
dP
dV
EFL
efl
ENDFILE
EVAL
expression1
expression2
expression3
FNCLEVEL
FRETURN
freturn
gcd
getobj
gimpel
griswold
i,j
i,k
k,j
kernighan
knuth
LE
lseek
Macrospitbol
MAXLNGTH
namemap
nobj
NOTANY
NRETURN
nreturn
obj
optblanks
P1&&P2
P1a
poage
POS
pre
proc1
proc1.h
proc2
proc2.h
qel
ratfor
ratsno
REM
rem.q
ritchie
RPOS
RTAB
sliteral
SNOBOL4
snobol4
Snocone
snocone
Snocone's
spitbol
square.end
statement1
statement2
STCOUNT
STLIMIT
struct
suc
term,1000
th
thompson
tl
unix
unqalphabet
usr
volume1
Yacc
zeroes
