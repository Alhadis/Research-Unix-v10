0,ta
0,tb
a,b
A.c
A.end
A.ne
A.nw
A.s
A.se
A.start
A.sw
a.tl
A:arc
a:arrow
A:circle
A:rect
acm
axx
axy
B.c
B.n
b.tl
b:arrow
bht
bot
bp
bro
bro.nw
bro.sw
bro:rect
btree
bu
bwd
c1,p1
c1,p1,p2,p3,p4,p5,r1,tp,bp,ta,tb
cis
colwid
conj
cstr
DV
e.g
eldest.nw
eldest.sw
eldest:rect
EQ
EQN
eqn
first.e
first.ht
first.info.hook
first.info.sw,first.next.se
first.ne
first.ne,first.se
first.next
first.next.c
first.next.ne,first.next.se
first.se
first.sw,first.se
first.w
gridline
gsize
hd
headang
headvec
hmv
ht
ibfile
id
idth
IE
im
info.nw
info.se
info.sw
int
inth
inth.e
inth.w,inth.e
inx
iny
ipth
ipth.e
ipth.w
isoceles
ith
ith.e
knuth
last.info.hook
last.info.sw
last.sw
last.w
leftpt
lesk
lht
libfile
listnode
llength
loc
lwd
Mashey
maxx
maxy
METAFONT
metafont
midang
midd
miny
ne
neg
new.info.hook
new.info.nw
new.next
new.next.c
new.nw
new.w
next.ne
next.nw
next.se
next.sw
next:rect
noerase
nw
nw,ne
obbox
olwid
opaqued
opaqueing
Opaquing
opaquing
pavlidis
perp
PIC
pic
poly
pos
PS
ps
pt1
pt2
pt3
pt4
pt5
r.c
r.e
r.s
r.w
radius,radius
rect
rh
rightpt
root.ne
root.nw
root.nw,root.sw
root.se
root.sw
root.sw,root.se
root:rect
rw
se
second.e
second.w,second.e
start,end
startang
sw
sw,se
T.z1
T.z2
T.z3
ta
tb
TBL
tbl
tf
tl
top,bot
tp
var
vert
vmv
VS
wd
wyk
yeserase
youngest.nw
youngest.se
youngest.sw
youngest:rect
ZAP.center
ZAP:circle
